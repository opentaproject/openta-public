Välkommen till uppgiftssystemet för {{course_name}}!

Ditt konto har användarnamn {{ username }} men är inte aktiverat än. Använd länken nedan för att aktivera och välja lösenord.
{{ activate_url }}

Efter aktivering kommer du automatiskt till inloggning som du senare hittar på adressen
{{ course_url }}

Om det uppstår frågor eller problem kan du svara på detta mail.

Lycka till!

Ps. Systemet är under aktiv utveckling, om du har synpunkter eller förslag på förbättringar får du gärna höra av dig.
